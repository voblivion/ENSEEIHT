library IEEE;
library UNISIM;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity clock28 is
	port (
		rst : in std_logic ;
		clk : in std_logic ;
		s : out std_logic_vector (27 downto 0)
	);
end clock28;

architecture synthesis of clock28 is

	-- submodules declarations
	component clock4
		port (
			rst : in std_logic ;
			clk : in std_logic ;
			s : out std_logic_vector (3 downto 0)
		) ;
	end component ;

	-- buffer signals declarations
	signal s_int : std_logic_vector (27 downto 0) ;

	-- internal signals declarations
	signal n3 : std_logic ;
	signal n7 : std_logic ;
	signal n11 : std_logic ;
	signal n15 : std_logic ;
	signal n19 : std_logic ;
	signal n23 : std_logic ;

begin

	-- buffer signals assignations
	s(27 downto 0) <= s_int(27 downto 0) ;

	-- concurrent statements
	n3 <= not s_int(3) ;
	n7 <= not s_int(7) ;
	n11 <= not s_int(11) ;
	n15 <= not s_int(15) ;
	n19 <= not s_int(19) ;
	n23 <= not s_int(23) ;

	-- components instanciations
	clock4_0 : clock4 port map (rst, clk, s_int(3 downto 0)) ;
	clock4_1 : clock4 port map (rst, n3, s_int(7 downto 4)) ;
	clock4_2 : clock4 port map (rst, n7, s_int(11 downto 8)) ;
	clock4_3 : clock4 port map (rst, n11, s_int(15 downto 12)) ;
	clock4_4 : clock4 port map (rst, n15, s_int(19 downto 16)) ;
	clock4_5 : clock4 port map (rst, n19, s_int(23 downto 20)) ;
	clock4_6 : clock4 port map (rst, n23, s_int(27 downto 24)) ;

end synthesis;
