library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity addbin_comm is
    port (
        mclk : in std_logic ;
        pdb : inout std_logic_vector (7 downto 0) ;
        astb : in std_logic ;
        dstb : in std_logic ;
        pwr : in std_logic ;
        pwait : out std_logic;
        btn : in std_logic_vector (1 downto 0) ;

        sw : in std_logic_vector (7 downto 7)

) ;
end addbin_comm ;

architecture synthesis of addbin_comm is

    -- submodules declarations
    component commUSB
        port (
            mclk     : in std_logic;
            pdb      : inout std_logic_vector(7 downto 0);
            astb     : in std_logic;
            dstb     : in std_logic;
            pwr      : in std_logic;
            pwait    : out std_logic;
            pc2board : out std_logic_vector(127 downto 0);
            board2pc : in std_logic_vector(127 downto 0)
        ) ;
    end component ;
	component addbin
		port (
			btn : in std_logic_vector (1 downto 0) ;
			sw : in std_logic_vector (7 downto 7) ;
			s : out std_logic ;
			cout : out std_logic
		) ;
	end component ;

    -- internal signals declarations
    signal pc2board : std_logic_vector (127 downto 0) ;
    signal board2pc : std_logic_vector (127 downto 0) ;
    signal s : std_logic ;
    signal cout : std_logic ;

begin

    -- combinatorial statements
    board2pc(0) <= s ;
    board2pc(1) <= cout ;

    -- components instanciations
    commUSB_0 : commUSB port map (mclk, pdb(7 downto 0), astb, dstb, pwr, pwait, pc2board(127 downto 0), board2pc(127 downto 0)) ;
    addbin_0 : addbin port map (btn(1 downto 0), sw(7 downto 7), s, cout) ;


end synthesis;
